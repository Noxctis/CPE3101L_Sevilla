// ======================================================================
// File:          Adder4bit.v
// Author:        Chrys Sean T. Sevilla
// Class:         CPE 3101L
// Group/Sched:   Group 4 Fri 10:30 - 1:30 PM
// Description:   Structural 4-bit ripple-carry adder using FullAdder cells
// ======================================================================

`timescale 1 ns / 1 ps

// ---------------------- Half Adder (gate primitives) -------------------
module HalfAdder (x, y, C, S);
  input  x, y;
  output C, S;

  xor X1 (S, x, y);
  and A1 (C, x, y);
endmodule

// ------------------------ Full Adder (structural) ----------------------
module FullAdder (Cin, A, B, FaS, FaC);
  input  Cin, A, B;
  output FaS, FaC;
  wire   C1, S1, C2;

  // First half adder: adds A and B
  HalfAdder HA1 (A, B, C1, S1);

  // Second half adder: adds S1 and Cin
  HalfAdder HA2 (S1, Cin, C2, FaS);

  // Final carry output
  or O1 (FaC, C1, C2);
endmodule

// --------------------------- 4-bit Adder -------------------------------
// Ripple-carry adder using four FullAdder instances
module Adder4Bit (A, B, C_in, S, C_out);
  input  [3:0] A, B;  // Unsigned preferred in waveform view
  input        C_in;
  output [3:0] S;
  output       C_out;

  wire C1, C2, C3;

  // LSB to MSB ripple
  FullAdder FA0 (C_in, A[0], B[0], S[0], C1);
  FullAdder FA1 (C1,   A[1], B[1], S[1], C2);
  FullAdder FA2 (C2,   A[2], B[2], S[2], C3);
  FullAdder FA3 (C3,   A[3], B[3], S[3], C_out);
endmodule
