module ClockDivider (
    input wire clk_in,      // 50 MHz input clock
    input wire nReset,      // Active-low asynchronous reset
    output reg clk_out      // Divided clock output
);

    // Calculate division factor:
    // 50 MHz / 2 Hz = 25,000,000 cycles per half-period
    parameter DIV_FACTOR = 25_000_000; // For FPGA
    // For simulation, use smaller value like 10 or 20

    reg [24:0] counter; // Enough bits for 25 million

    always @(posedge clk_in or negedge nReset) begin
        if (!nReset) begin
            counter <= 0;
            clk_out <= 0;
        end else begin
            if (counter == DIV_FACTOR - 1) begin
                counter <= 0;
                clk_out <= ~clk_out; // Toggle output
            end else begin
                counter <= counter + 1;
            end
        end
    end

endmodule
