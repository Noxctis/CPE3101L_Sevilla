module tb_ClockDivider;

    reg clk_in, nReset;
    wire clk_out;

    // Instantiate Clock Divider with smaller factor for simulation
    ClockDivider #(.DIV_FACTOR(10)) uut (
        .clk_in(clk_in),
        .nReset(nReset),
        .clk_out(clk_out)
    );

    // Generate input clock (simulate 50 MHz scaled down)
    initial begin
        clk_in = 0;
        forever #1 clk_in = ~clk_in; // 1 time unit period
    end

    initial begin
        $display("Time\tclk_in\tnReset\tclk_out");
        $monitor("%0t\t%b\t%b\t%b", $time, clk_in, nReset, clk_out);

        // Assert reset
        nReset = 0; #5;
        nReset = 1;

        // Let clock run for a while
        #200;

        $stop;
    end

endmodule