/*
File:					tb_HalfAdder.v
Author:				Chrys Sean T. Sevilla
Class:				CPE 3101L
Group/Schedule: 	Group 4 Fri 10:30 - 1:30 PM
Description:		Testbench file for HalfAdderAdder.v

*/

`timescale 1 ns/ 1ps

module tb_HalfAdder();

	reg	x, y;
	wire	C, S;
	
	HalfAdder UUT (x,y,C,S);
	
	initial
	begin
		x = 0;	y = 0;	#10
		x = 0;	y = 1;	#10
		x = 1;	y = 0;	#10
		x = 1;	y = 1;	#50
		
		$stop;
	end
	
endmodule